// define this macro to enable fast behavior simulation
// for flash by skipping SPI transfers
// `define FAST_FLASH

module spi_top_apb #(
    parameter flash_addr_start = 32'h30000000,
    parameter flash_addr_end   = 32'h3fffffff,
    parameter spi_ss_num       = 8
) (
    input         clock,
    input         reset,
    input  [31:0] in_paddr,
    input         in_psel,
    input         in_penable,
    input  [ 2:0] in_pprot,
    input         in_pwrite,
    input  [31:0] in_pwdata,
    input  [ 3:0] in_pstrb,
    output        in_pready,
    output [31:0] in_prdata,
    output        in_pslverr,

    output                  spi_sck,
    output [spi_ss_num-1:0] spi_ss,
    output                  spi_mosi,
    input                   spi_miso,
    output                  spi_irq_out
);

`ifdef FAST_FLASH

  wire [31:0] data;
  parameter invalid_cmd = 8'h0;
  flash_cmd flash_cmd_i (
      .clock(clock),
      .valid(in_psel && !in_penable),
      .cmd  (in_pwrite ? invalid_cmd : 8'h03),
      .addr ({8'b0, in_paddr[23:2], 2'b0}),
      .data (data)
  );
  assign spi_sck     = 1'b0;
  assign spi_ss      = 8'b0;
  assign spi_mosi    = 1'b1;
  assign spi_irq_out = 1'b0;
  assign in_pslverr  = 1'b0;
  assign in_pready   = in_penable && in_psel && !in_pwrite;
  assign in_prdata   = data[31:0];

`else

  spi_top u0_spi_top (
      .wb_clk_i(clock),
      .wb_rst_i(reset),
      .wb_adr_i(in_paddr[4:0]),
      .wb_dat_i(in_pwdata),
      .wb_dat_o(in_prdata),
      .wb_sel_i(in_pstrb),
      .wb_we_i (in_pwrite),
      .wb_stb_i(in_psel),
      .wb_cyc_i(in_penable),
      .wb_ack_o(in_pready),
      .wb_err_o(in_pslverr),
      .wb_int_o(spi_irq_out),

      .ss_pad_o  (spi_ss),
      .sclk_pad_o(spi_sck),
      .mosi_pad_o(spi_mosi),
      .miso_pad_i(spi_miso)
  );

`endif  // FAST_FLASH

endmodule
